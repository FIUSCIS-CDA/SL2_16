///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SPLICE_SL2
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A (16-bit)
reg[15:0] A;
///////////////////////////////////////////////////////////////////////////////////
// Output: S (18-bit)
wire[17:0] S;
///////////////////////////////////////////////////////////////////////////////////

SPLICE_SL2 mySL2(.A(A), .Y(S));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: A=3782
$display("Test: A=3782");
A=3782;   #10; 
verifyEqual32(S, A*4);
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule