///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SL2_16
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A (16-bit)
reg[15:0] A;
///////////////////////////////////////////////////////////////////////////////////
// Output: Y (18-bit)
wire[17:0] Y;
///////////////////////////////////////////////////////////////////////////////////

SL2_16 mySL2(.A(A), .Y(Y));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: A=3782
$display("Test: A=3782");
A=3782;   #10; 
verifyEqual32(Y, A*4);
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule
